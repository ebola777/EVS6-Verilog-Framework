///////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer: Shawn Chang (ebola777@yahoo.com.tw)
//
// Create Date: 20:01:00 04/07/2015
// Design Name:
// Module Name:
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////
`ifndef _characters_vh_
`define _characters_vh_

// Used to suppress unused leftmost bit of 8-bit ASCII characters.
`define CHAR_FILLED 8'b1111_1110
`define CHAR_SPACE 8'b1111_1111

`endif
