///////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer: Shawn Chang (ebola777@yahoo.com.tw)
//
// Create Date: 20:01:00 04/07/2015
// Design Name:
// Module Name:
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////
`ifndef _directives_vh_
`define _directives_vh_

`include "frequency.vh"
`include "io.vh"
`include "lcd.vh"
`include "audio.vh"
`include "debounce.vh"
`include "data_type.vh"
`include "characters.vh"

`endif
