///////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer: Shawn Chang (ebola777@yahoo.com.tw)
//
// Create Date: 20:01:00 04/07/2015
// Design Name:
// Module Name:
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////
`ifndef _audio_vh_
`define _audio_vh_

`define AUDIO_BIT_DEPTH 3
`define AUDIO_BIT_WIDTH_DATA 8

`define AUDIO_INITIAL_VOLUME 6'b00_0000

`endif
