///////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer: Shawn Chang (ebola777@yahoo.com.tw)
//
// Create Date: 20:01:00 04/07/2015
// Design Name:
// Module Name:
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////
`ifndef _debounce_vh_
`define _debounce_vh_

`define DEBOUNCE_LENGTH_PUSHBUTTON 6
`define DEBOUNCE_LENGTH_PUSHBUTTON_BIT_WIDTH 3

`define DEBOUNCE_LENGTH_KEYBOARD 6
`define DEBOUNCE_LENGTH_KEYBOARD_BIT_WIDTH 3

`endif
